LIBRARY IEEE;
USE  IEEE.STD_LOGIC_1164.all;
USE  IEEE.STD_LOGIC_UNSIGNED.all;

ENTITY contador_2seg_vhdl IS
	PORT(clock,enable,reset : IN STD_LOGIC;
		 dos_seg : OUT STD_LOGIC;
		 Q : Buffer STD_LOGIC_VECTOR (1 downto 0));
END contador_2seg_vhdl;

ARCHITECTURE sol OF contador_2seg_vhdl IS
BEGIN

	PROCESS(clock,reset)
	BEGIN
		if reset='0' then Q<="00";dos_seg<='0';
  		elsif (clock'event and clock='1') then
			if enable='1' then
				if (Q="10") then Q<="00";dos_seg<='1';
				else Q<=Q+1;dos_seg<='0';
				end if;
			end if;
		end if;
	END PROCESS;
END sol;