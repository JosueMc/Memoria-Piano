LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;
USE IEEE.STD_LOGIC_ARITH.all;
USE IEEE.STD_LOGIC_UNSIGNED.all;


entity musicasave is
	port(modo: in std_logic_vector(4 downto 0);
	q0,q1,q2,q3,q4,q5,q6,q7,q8,q9: out std_logic_vector(6 downto 0));
end musicasave;
architecture sol of musicasave is
begin
		process(modo)
			begin
				if modo="00000" then --musica 0
					q0<="0000001";q1<="0000010";
					q2<="0000100";q3<="0001000";
					q4<="0010000";q5<="0100000";
					q6<="1000000";q7<="0000001";
					q8<="0000001";q9<="0000001";
				elsif modo="00001" then --musica 1
					q0<="0010000";q1<="0000010";
					q2<="0000010";q3<="0001000";
					q4<="0100000";q5<="0100000";
					q6<="0001000";q7<="0000001";
					q8<="0000100";q9<="1000000";
				elsif modo="00010" then --musica 2
					q0<="0000001";q1<="0000010";
					q2<="0010000";q3<="1000000";
					q4<="1000000";q5<="0001000";
					q6<="0001000";q7<="0100000";
					q8<="0000001";q9<="0000010";
				elsif modo="00011" then --musica 3
					q0<="0000001";q1<="0000010";
					q2<="0100000";q3<="0010000";
					q4<="1000000";q5<="0100000";
					q6<="0000001";q7<="0001000";
					q8<="0000001";q9<="0000100";
				elsif modo="00100" then --musica 4
					q0<="0010000";q1<="0001000";
					q2<="0000010";q3<="0001000";
					q4<="1000000";q5<="0100000";
					q6<="0000010";q7<="0001000";
					q8<="0100000";q9<="0010000";
				elsif modo="00101" then --musica 5
					q0<="0001000";q1<="0010000";
					q2<="0000100";q3<="0001000";
					q4<="0000100";q5<="0100000";
					q6<="0001000";q7<="1000000";
					q8<="0000001";q9<="0000010";
				elsif modo="00110" then --musica 6
					q0<="0000010";q1<="0000100";
					q2<="0000100";q3<="0010000";
					q4<="0010000";q5<="0100000";
					q6<="0001000";q7<="1000000";
					q8<="0000001";q9<="0000010";
				elsif modo="00111" then --musica 7
					q0<="0000100";q1<="0000001";
					q2<="0000100";q3<="0001000";
					q4<="0010000";q5<="0100000";
					q6<="1000000";q7<="0001000";
					q8<="0000001";q9<="0010000";
				elsif modo="01000" then --musica 8
					q0<="1000000";q1<="0000010";
					q2<="0000100";q3<="0001000";
					q4<="0010000";q5<="0100000";
					q6<="1000000";q7<="0000001";
					q8<="0000001";q9<="1000000";
				elsif modo="01001" then --musica 9
					q0<="1000000";q1<="0001000";
					q2<="0000100";q3<="0001000";
					q4<="0010000";q5<="0100000";
					q6<="1000000";q7<="1000000";
					q8<="0001000";q9<="0000001";
				elsif modo="01010" then --musica 10
					q0<="1000000";q1<="0000010";
					q2<="0000100";q3<="0001000";
					q4<="0010000";q5<="0100000";
					q6<="1000000";q7<="0000001";
					q8<="0000001";q9<="0100000";
				elsif modo="01011" then --musica 11
					q0<="0000100";q1<="1000000";
					q2<="0000100";q3<="0001000";
					q4<="1000000";q5<="0100000";
					q6<="1000000";q7<="0000010";
					q8<="0000001";q9<="0100000";
				elsif modo="01100" then --musica 12
					q0<="0000001";q1<="0100000";
					q2<="0000010";q3<="0001000";
					q4<="0010000";q5<="0100000";
					q6<="0000010";q7<="0000001";
					q8<="0000010";q9<="0000001";
				elsif modo="01101" then --musica 13
					q0<="0000001";q1<="1000000";
					q2<="0000100";q3<="0001000";
					q4<="1000000";q5<="0100000";
					q6<="1000000";q7<="1000000";
					q8<="0000001";q9<="1000000";
				elsif modo="01110" then --musica 14
					q0<="0000001";q1<="0000010";
					q2<="0000100";q3<="0001000";
					q4<="0010000";q5<="0100000";
					q6<="1000000";q7<="0000001";
					q8<="0000001";q9<="0000001";
				elsif modo="01111" then --musica 15
					q0<="0000001";q1<="1000000";
					q2<="0000100";q3<="1000000";
					q4<="0010000";q5<="0000100";
					q6<="1000000";q7<="0000001";
					q8<="0000001";q9<="0000100";
				elsif modo="10000" then --musica 16
					q0<="0000001";q1<="0000010";
					q2<="0000100";q3<="0000001";
					q4<="0010000";q5<="0100000";
					q6<="1000000";q7<="0000001";
					q8<="0000001";q9<="1000000";
				elsif modo="10001" then --musica 17
					q0<="0000001";q1<="0000010";
					q2<="0000100";q3<="0001000";
					q4<="0010000";q5<="0100000";
					q6<="1000000";q7<="0000001";
					q8<="0000001";q9<="0000001";
				elsif modo="10010" then --musica 18
					q0<="0000010";q1<="0000010";
					q2<="0000100";q3<="0001000";
					q4<="0010000";q5<="0000100";
					q6<="0000010";q7<="0000001";
					q8<="0000001";q9<="0000010";
				elsif modo="10011" then --musica 19
					q0<="0000001";q1<="0000010";
					q2<="0000100";q3<="0001000";
					q4<="0010000";q5<="0100000";
					q6<="1000000";q7<="0010000";
					q8<="0000100";q9<="0000001";
				end if;
	end process;
end sol;